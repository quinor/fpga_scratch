`timescale 1ns / 1ps

module vga(
    input clk,
    output [3:0] vgaRed, // delayed by 2
    output [3:0] vgaGreen, // delatyed by 2
    output [3:0] vgaBlue, // delayed by 2
    output Vsync, // delayed by 2
    output Hsync, // delayed by 2
    input write_clk,
    input [7:0] write_posx,
    input [5:0] write_posy,
    input [31:0] write_value,
    input write_enable,
    input [5:0] v_offset
    );

localparam W = 1280;
localparam HFRONT = 72;
localparam HSYNC = 80;
localparam HBACK = 216;
localparam LINE = W + HFRONT + HSYNC + HBACK;

localparam H = 720;
localparam VFRONT = 3;
localparam VSYNC = 5;
localparam VBACK = 22;
localparam PAGE = H + VFRONT + VSYNC + VBACK;


wire vga_clk;
wire feedback;

PLLE2_BASE #(
    .CLKFBOUT_MULT(52), // Multiply value for all CLKOUT, (2-64)
    .CLKIN1_PERIOD(10.0), // Input clock period in ns to ps resolution (i.e. 33.333 is 30 MHz).
    .CLKOUT0_DIVIDE(14),
    .DIVCLK_DIVIDE(5),
    .STARTUP_WAIT("TRUE") // Delay DONE until PLL Locks, ("TRUE"/"FALSE")
) PLLE2_BASE_inst (
    .CLKOUT0(vga_clk), // 1-bit output: CLKOUT0
    .CLKFBOUT(feedback), // 1-bit output: Feedback clock
    .CLKIN1(clk), // 1-bit input: Input clock
    .CLKFBIN(feedback) // 1-bit input: Feedback clock
);


wire [11:0] index_addr; // delayed by 1
wire [7:0] index_value; // delayed by 2

BRAM_SDP_MACRO #(
    .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb"
    .DEVICE("7SERIES"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6", "7SERIES"
    .WRITE_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
    .READ_WIDTH(8), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
    .INIT_00(256'h000000007e818199bd8181a5817e000000000000000000000000000000000000),
    .INIT_01(256'h00000000081c3e7f7f7f7f3600000000000000007effffe7c3ffffdbff7e0000),
    .INIT_02(256'h000000003c1818e7e7e73c3c180000000000000000081c3e7f3e1c0800000000),
    .INIT_03(256'h000000000000183c3c18000000000000000000003c18187effff7e3c18000000),
    .INIT_04(256'h00000000003c664242663c0000000000ffffffffffffe7c3c3e7ffffffffffff),
    .INIT_05(256'h000000001e333333331e4c5870780000ffffffffffc399bdbd99c3ffffffffff),
    .INIT_06(256'h00000000070f0e0c0c0c0cfcccfc00000000000018187e183c666666663c0000),
    .INIT_07(256'h000000001818db3ce73cdb18180000000000000367e7e6c6c6c6c6fec6fe0000),
    .INIT_08(256'h00000000406070787c7f7c7870604000000000000103070f1f7f1f0f07030100),
    .INIT_09(256'h000000006666006666666666666600000000000000183c7e1818187e3c180000),
    .INIT_0A(256'h0000003e63301c366363361c06633e0000000000d8d8d8d8d8dedbdbdbfe0000),
    .INIT_0B(256'h000000007e183c7e1818187e3c180000000000007f7f7f7f0000000000000000),
    .INIT_0C(256'h00000000183c7e18181818181818000000000000181818181818187e3c180000),
    .INIT_0D(256'h0000000000000c067f060c000000000000000000000018307f30180000000000),
    .INIT_0E(256'h00000000000014367f361400000000000000000000007f030303000000000000),
    .INIT_0F(256'h0000000000081c1c3e3e7f7f0000000000000000007f7f3e3e1c1c0800000000),
    .INIT_10(256'h000000001818001818183c3c3c18000000000000000000000000000000000000),
    .INIT_11(256'h0000000036367f3636367f363600000000000000000000000000002466666600),
    .INIT_12(256'h000000006163060c1830634300000000000018183e636160603e0343633e1818),
    .INIT_13(256'h0000000000000000000000060c0c0c00000000006e3333333b6e1c36361c0000),
    .INIT_14(256'h000000000c18303030303030180c00000000000030180c0c0c0c0c0c18300000),
    .INIT_15(256'h00000000000018187e18180000000000000000000000663cff3c660000000000),
    .INIT_16(256'h00000000000000007f000000000000000000000c181818000000000000000000),
    .INIT_17(256'h000000000103060c183060400000000000000000181800000000000000000000),
    .INIT_18(256'h000000007e1818181818181e1c180000000000001c3663636b6b6363361c0000),
    .INIT_19(256'h000000003e636060603c6060633e0000000000007f6303060c183060633e0000),
    .INIT_1A(256'h000000003e636060603f0303037f000000000000783030307f33363c38300000),
    .INIT_1B(256'h000000000c0c0c0c18306060637f0000000000003e636363633f0303061c0000),
    .INIT_1C(256'h000000001e306060607e6363633e0000000000003e636363633e6363633e0000),
    .INIT_1D(256'h000000000c181800000018180000000000000000001818000000181800000000),
    .INIT_1E(256'h000000000000007e00007e0000000000000000006030180c060c183060000000),
    .INIT_1F(256'h000000001818001818183063633e000000000000060c18306030180c06000000),
    .INIT_20(256'h00000000636363637f6363361c080000000000003e033b7b7b7b63633e000000),
    .INIT_21(256'h000000003c66430303030343663c0000000000003f666666663e6666663f0000),
    .INIT_22(256'h000000007f664606161e1646667f0000000000001f36666666666666361f0000),
    .INIT_23(256'h000000005c6663637b030343663c0000000000000f060606161e1646667f0000),
    .INIT_24(256'h000000003c18181818181818183c00000000000063636363637f636363630000),
    .INIT_25(256'h00000000676666361e1e366666670000000000001e3333333030303030780000),
    .INIT_26(256'h0000000063636363636b7f7f77630000000000007f66460606060606060f0000),
    .INIT_27(256'h000000003e63636363636363633e00000000000063636363737b7f6f67630000),
    .INIT_28(256'h000070303e7b6b6363636363633e0000000000000f060606063e6666663f0000),
    .INIT_29(256'h000000003e636360301c0663633e00000000000067666666363e6666663f0000),
    .INIT_2A(256'h000000003e6363636363636363630000000000003c1818181818185a7e7e0000),
    .INIT_2B(256'h0000000036777f6b6b6b63636363000000000000081c36636363636363630000),
    .INIT_2C(256'h000000003c181818183c666666660000000000006363363e1c1c3e3663630000),
    .INIT_2D(256'h000000003c0c0c0c0c0c0c0c0c3c0000000000007f6343060c183061637f0000),
    .INIT_2E(256'h000000003c30303030303030303c000000000000406070381c0e070301000000),
    .INIT_2F(256'h0000ff0000000000000000000000000000000000000000000000000063361c08),
    .INIT_30(256'h000000006e3333333e301e000000000000000000000000000000000030180c00),
    .INIT_31(256'h000000003e63030303633e0000000000000000003e66666666361e0606070000),
    .INIT_32(256'h000000003e6303037f633e0000000000000000006e33333333363c3030380000),
    .INIT_33(256'h001e33303e33333333336e0000000000000000001e0c0c0c0c1e0c4c6c380000),
    .INIT_34(256'h000000003c18181818181c00181800000000000067666666666e360606070000),
    .INIT_35(256'h000000006766361e1e36660606070000003c6666606060606060700060600000),
    .INIT_36(256'h00000000636b6b6b6b7f370000000000000000003c18181818181818181c0000),
    .INIT_37(256'h000000003e63636363633e0000000000000000006666666666663b0000000000),
    .INIT_38(256'h007830303e33333333336e0000000000000f06063e66666666663b0000000000),
    .INIT_39(256'h000000003e63301c06633e0000000000000000000f060606666e3b0000000000),
    .INIT_3A(256'h000000006e333333333333000000000000000000386c0c0c0c0c3f0c0c080000),
    .INIT_3B(256'h00000000367f6b6b6b63630000000000000000001c3663636363630000000000),
    .INIT_3C(256'h001f30607e63636363636300000000000000000063361c1c1c36630000000000),
    .INIT_3D(256'h0000000070181818180e181818700000000000007f63060c18337f0000000000),
    .INIT_3E(256'h000000000e18181818701818180e000000000000181818181818181818180000),
    .INIT_3F(256'h00000000007f636363361c0800000000000000000000000000000000003b6e00),
    .INIT_40(256'h000000006e333333333333000033000000000e183c66430303030343663c0000),
    .INIT_41(256'h000000006e3333333e301e00361c0800000000003e6303037f633e000c183000),
    .INIT_42(256'h000000006e3333333e301e00180c0600000000006e3333333e301e0000330000),
    .INIT_43(256'h00000e183e63030303633e0000000000000000006e3333333e301e001c361c00),
    .INIT_44(256'h000000003e6303037f633e0000630000000000003e6303037f633e00361c0800),
    .INIT_45(256'h000000003c18181818181c0000660000000000003e6303037f633e00180c0600),
    .INIT_46(256'h000000003c18181818181c00180c0600000000003c18181818181c00663c1800),
    .INIT_47(256'h00000000636363637f63361c081c361c000000006363637f6363361c08006300),
    .INIT_48(256'h00000000761b1b7e6c6c370000000000000000007f6646161e1646667f001830),
    .INIT_49(256'h000000003e63636363633e00361c08000000000073333333337f3333367c0000),
    .INIT_4A(256'h000000003e63636363633e00180c0600000000003e63636363633e0000630000),
    .INIT_4B(256'h000000006e33333333333300180c0600000000006e33333333333300331e0c00),
    .INIT_4C(256'h000000003e636363636363633e006300001e30607e6363636363630000630000),
    .INIT_4D(256'h0000000018183e63030303633e181800000000003e6363636363636363006300),
    .INIT_4E(256'h000000001818187e187e183c66660000000000003f67060606060f0626361c00),
    .INIT_4F(256'h000000000e1b1818187e181818d8700000000000633333337b33231f33331f00),
    .INIT_50(256'h000000003c18181818181c000c183000000000006e3333333e301e00060c1800),
    .INIT_51(256'h000000006e33333333333300060c1800000000003e63636363633e00060c1800),
    .INIT_52(256'h00000000636363737b7f6f6763003b6e000000006666666666663b003b6e0000),
    .INIT_53(256'h00000000000000003e001c36361c000000000000000000007e007c36363c0000),
    .INIT_54(256'h0000000000030303037f000000000000000000003e636303060c0c000c0c0000),
    .INIT_55(256'h00007c1830613b060c183666460706000000000000606060607f000000000000),
    .INIT_56(256'h00000000183c3c3c181818001818000000006060fc5973660c18366646070600),
    .INIT_57(256'h0000000000001b366c361b00000000000000000000006c361b366c0000000000),
    .INIT_58(256'h55aa55aa55aa55aa55aa55aa55aa55aa22882288228822882288228822882288),
    .INIT_59(256'h18181818181818181818181818181818eebbeebbeebbeebbeebbeebbeebbeebb),
    .INIT_5A(256'h18181818181818181f181f181818181818181818181818181f18181818181818),
    .INIT_5B(256'h6c6c6c6c6c6c6c6c7f000000000000006c6c6c6c6c6c6c6c6f6c6c6c6c6c6c6c),
    .INIT_5C(256'h6c6c6c6c6c6c6c6c6f606f6c6c6c6c6c18181818181818181f181f0000000000),
    .INIT_5D(256'h6c6c6c6c6c6c6c6c6f607f00000000006c6c6c6c6c6c6c6c6c6c6c6c6c6c6c6c),
    .INIT_5E(256'h00000000000000007f6c6c6c6c6c6c6c00000000000000007f606f6c6c6c6c6c),
    .INIT_5F(256'h18181818181818181f0000000000000000000000000000001f181f1818181818),
    .INIT_60(256'h0000000000000000ff181818181818180000000000000000f818181818181818),
    .INIT_61(256'h1818181818181818f8181818181818181818181818181818ff00000000000000),
    .INIT_62(256'h1818181818181818ff181818181818180000000000000000ff00000000000000),
    .INIT_63(256'h6c6c6c6c6c6c6c6cec6c6c6c6c6c6c6c1818181818181818f818f81818181818),
    .INIT_64(256'h6c6c6c6c6c6c6c6cec0cfc00000000000000000000000000fc0cec6c6c6c6c6c),
    .INIT_65(256'h6c6c6c6c6c6c6c6cef00ff00000000000000000000000000ff00ef6c6c6c6c6c),
    .INIT_66(256'h0000000000000000ff00ff00000000006c6c6c6c6c6c6c6cec0cec6c6c6c6c6c),
    .INIT_67(256'h0000000000000000ff00ff18181818186c6c6c6c6c6c6c6cef00ef6c6c6c6c6c),
    .INIT_68(256'h1818181818181818ff00ff00000000000000000000000000ff6c6c6c6c6c6c6c),
    .INIT_69(256'h0000000000000000fc6c6c6c6c6c6c6c6c6c6c6c6c6c6c6cff00000000000000),
    .INIT_6A(256'h1818181818181818f818f800000000000000000000000000f818f81818181818),
    .INIT_6B(256'h6c6c6c6c6c6c6c6cff6c6c6c6c6c6c6c6c6c6c6c6c6c6c6cfc00000000000000),
    .INIT_6C(256'h00000000000000001f181818181818181818181818181818ff18ff1818181818),
    .INIT_6D(256'hffffffffffffffffffffffffffffffff1818181818181818f800000000000000),
    .INIT_6E(256'h0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0fffffffffffffffffff00000000000000),
    .INIT_6F(256'h000000000000000000fffffffffffffff0f0f0f0f0f0f0f0f0f0f0f0f0f0f0f0),
    .INIT_70(256'h0000000033636363331b3333331e0000000000006e3b1b1b1b3b6e0000000000),
    .INIT_71(256'h000000003636363636367f0000000000000000000303030303030363637f0000),
    .INIT_72(256'h000000000e1b1b1b1b1b7e0000000000000000007f63060c18180c06637f0000),
    .INIT_73(256'h000000001818181818183b6e00000000000306063e6666666666660000000000),
    .INIT_74(256'h000000001c366363637f6363361c0000000000007e183c666666663c187e0000),
    .INIT_75(256'h000000003c666666667c30180c780000000000007736363636636363361c0000),
    .INIT_76(256'h0000000003067ecfdbdb7e60c00000000000000000007edbdbdb7e0000000000),
    .INIT_77(256'h0000000063636363636363633e00000000000000380c0606063e06060c380000),
    .INIT_78(256'h000000007e000018187e18180000000000000000007f00007f00007f00000000),
    .INIT_79(256'h000000007e0030180c060c1830000000000000007e000c18306030180c000000),
    .INIT_7A(256'h0000000e1b1b1b1818181818181818181818181818181818181818d8d8700000),
    .INIT_7B(256'h0000000000003b6e003b6e000000000000000000000018007e00180000000000),
    .INIT_7C(256'h0000000000000018180000000000000000000000000000000000001c36361c00),
    .INIT_7D(256'h00000000383c3636373030303030f00000000000000000001800000000000000),
    .INIT_7E(256'h0000000000000000007e4c1830663c000000000000000000006c6c6c6c6c3600),
    .INIT_7F(256'h0000000000000000000000000000000000000000007e7e7e7e7e7e7e00000000),
    .WRITE_MODE("WRITE_FIRST") // Specify "READ_FIRST" for same clock or synchronous clocks
// Specify "WRITE_FIRST for asynchronous clocks on ports
) block1 (
    .DO(index_value), // Output read data port, width defined by READ_WIDTH parameter
    .RDADDR(index_addr), // Input read address, width defined by read port depth
    .RDCLK(vga_clk), // 1-bit input read clock
    .RDEN(1), // 1-bit input read port enable

    .RST(0), // 1-bit input reset

    .DI(0), // Input write data port, width defined by WRITE_WIDTH parameter
    .WE(0), // Input write enable, width defined by write port depth
    .WRADDR(0), // Input write address, width defined by write port depth
    .WRCLK(0), // 1-bit input write clock
    .WREN(0), // 1-bit input write port enable
    .REGCE(0)
);


wire [12:0] framebuffer_addr;
wire [31:0] framebuffer_value; // delayed by 1
wire [11:0] col1, col2; // delayed by 2

delay #(.BITS(24), .DELAY(1)) (vga_clk, {col1, col2}, framebuffer_value[31:8]);

wire [12:0] write_addr;

assign write_addr = write_posx + (write_posy << 7) + (write_posy << 5);

reg [31:0] write_value_1;
reg [12:0] write_addr_1;
reg write_enable_1;

always @(posedge write_clk) begin
    write_value_1 <= write_value;
    write_addr_1 <= write_addr;
    write_enable_1 <= write_enable;
end

blockram #(
    .WIDTH(2)
) br (
    vga_clk, framebuffer_addr, framebuffer_value,
    write_clk, write_addr_1, write_value_1, write_enable_1
);


reg [15:0] v_pos, h_pos;
wire [11:0] rgb;

wire display_enable; // delayed by 2

delay #(.BITS(1), .DELAY(2)) (vga_clk, Hsync, ~(h_pos >= W + HFRONT & h_pos < W + HFRONT + HSYNC));
delay #(.BITS(1), .DELAY(2)) (vga_clk, Vsync, ~(v_pos >= H + VFRONT & v_pos < H + VFRONT + VSYNC));
delay #(.BITS(1), .DELAY(2)) (vga_clk, display_enable, v_pos < H & h_pos < W);

assign {vgaRed, vgaGreen, vgaBlue} = display_enable ? rgb : 0;


(* ASYNC_REG = "TRUE" *) reg [5:0] off_sync_0, off_sync_1, off_sync_2, off_sync_3, off_sync_4;
reg [5:0] v_offset_current;

always @(posedge vga_clk) begin
    off_sync_0 <= v_offset;
    off_sync_1 <= off_sync_0;
    off_sync_2 <= off_sync_1;
    off_sync_3 <= off_sync_2;
    off_sync_4 <= off_sync_3;
    if (
        Vsync == 0
        && off_sync_0 == off_sync_1
        && off_sync_1 == off_sync_2
        && off_sync_2 == off_sync_3
        && off_sync_3 == off_sync_4
    )
        v_offset_current <= off_sync_4;
end


wire [12:0] v_pos_offset;

simplemod #(.BITS(13), .MOD(45)) mod (v_pos_offset, {1'b0, v_pos[15:4] + v_offset_current});

assign framebuffer_addr = h_pos[15:3] + (v_pos_offset << 7) + (v_pos_offset << 5);


wire [3:0] dy_d; // delayed by 1
wire [2:0] dx_d; // delayed by 2
delay #(.BITS(4), .DELAY(1)) (vga_clk, dy_d, v_pos[3:0]);
delay #(.BITS(3), .DELAY(2)) (vga_clk, dx_d, h_pos[2:0]);

assign index_addr = {framebuffer_value[7:0], dy_d};

assign rgb = index_value[dx_d] ? col1 : col2;

always @(posedge vga_clk) begin
    if (h_pos == LINE-1) begin
        h_pos <= 0;
        if (v_pos == PAGE-1)
            v_pos <= 0;
        else
            v_pos <= v_pos + 1;
    end else
        h_pos <= h_pos + 1;
end

endmodule
